/*

Copyright (c) 2014-2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`resetall
`timescale 1ns / 1ps
`default_nettype none

/*
 * FPGA top-level module
 */
module fpga (
    /*
     * Clock: 200MHz
     * Reset: Push button, active high
     */
    input  wire       clk_200mhz_p,
    input  wire       clk_200mhz_n,
    //input  wire       reset,

    /*
     * GPIO
     */
    input  wire       btnu,
    input  wire       btnl,
    input  wire       btnd,
    input  wire       btnr,
    input  wire       btnc,
    input  wire [3:0] sw,
    output wire [7:0] led,

    /*
     * Ethernet: 100BASE-T RMII
     */

    input  wire [1:0] phy_rxd,
    input  wire       phy_rx_er,
    input  wire       phy_crs_dv,
    output wire [1:0] phy_txd,
    output wire       phy_tx_en,
    output wire       phy_ref_clk,  //50Mhz reference clock
    output wire       phy_reset_n,
    inout  wire       rgmii_mdio_a,

    input  wire       macif_sel0,  

    /*
     * UART: 500000 bps, 8N1
     */
    input  wire       uart_rxd,
    output wire       uart_txd,
    output wire       uart_rts,
    input  wire       uart_cts
);
//tests
wire reset =  btnc;
wire phy_reset;
assign phy_reset_n = !phy_reset;
wire [7:0] led_out;
reg [26:0] clk_counter;
reg [26:0] clk_rx_counter;
reg clk_1Hz_rx;
reg clk_1Hz;

assign led[0] = 1'b0;
assign led[1] = 1'b1;
assign led[2] = reset;
assign led[3] = phy_reset_n;
assign led[4] = clk_1Hz;
assign led[5] = clk_1Hz_rx;
assign led[7:6] = led_out[7:6];


// Clock and reset
wire phy_int_n = 1'b0;
wire clk_200mhz_ibufg;

// Internal 125 MHz clock
wire clk_mmcm_out;
wire clk_int;
wire rst_int;

wire clk_200mhz_mmcm_out;
wire clk_200mhz_int;

// Reference clock for RMII
wire clk_50mhz_mmcm_out;
wire clk_50mhz_int;
wire phy_mii_tx_clk;

// Reference clock for MII
// wire clk_25mhz_mmcm_out;
// wire clk_25mhz_int;

wire mmcm_rst = reset;
wire mmcm_locked;
wire mmcm_clkfb;

assign phy_ref_clk = clk_50mhz_int;

//ila_0 
//RXPROBE(
//.clk(phy_rx_clk),
//.probe0(phy_rxd),
//.probe1(phy_rx_ctl)
//);



IBUFGDS
clk_200mhz_ibufgds_inst(
    .I(clk_200mhz_p),
    .IB(clk_200mhz_n),
    .O(clk_200mhz_ibufg)
);

//LUDO 1 Hz blink
always @(posedge clk_50mhz_int) begin
    if (clk_counter >= 50_000_000/2 - 1) begin
        clk_counter <= 0; // Reset counter when it reaches 
        clk_1Hz <= ~clk_1Hz;
    end else begin
        clk_counter <= clk_counter + 1; // Increment counter
    end
end
always @(posedge phy_mii_tx_clk) begin
    if (clk_rx_counter >= 25_000_000/2 - 1) begin
        clk_rx_counter <= 0; // Reset counter when it reaches
        clk_1Hz_rx <= ~clk_1Hz_rx;
    end else begin
        clk_rx_counter <= clk_rx_counter + 1; // Increment counter
    end
end


// MMCM instance
// 200 MHz in, 125 MHz out
// PFD range: 10 MHz to 500 MHz
// VCO range: 600 MHz to 1440 MHz
// M = 5, D = 1 sets Fvco = 1000 MHz (in range)
// Divide by 8 to get output frequency of 125 MHz
// Divide by 40 to get output frequency of 25 MHz
// Divide by 20 to get output frequency of 50 MHz
// Also need 200 MHz out for IODELAY
// 1000 / 5 = 200 MHz
MMCME2_BASE #(
    .BANDWIDTH("OPTIMIZED"),
    .CLKOUT0_DIVIDE_F(8),
    .CLKOUT0_DUTY_CYCLE(0.5),
    .CLKOUT0_PHASE(0),
    .CLKOUT1_DIVIDE(40),
    .CLKOUT1_DUTY_CYCLE(0.5),
    .CLKOUT1_PHASE(0),
    .CLKOUT2_DIVIDE(5),
    .CLKOUT2_DUTY_CYCLE(0.5),
    .CLKOUT2_PHASE(0),
    .CLKOUT3_DIVIDE(20),
    .CLKOUT3_DUTY_CYCLE(0.5),
    .CLKOUT3_PHASE(0),
    .CLKOUT4_DIVIDE(1),
    .CLKOUT4_DUTY_CYCLE(0.5),
    .CLKOUT4_PHASE(0),
    .CLKOUT5_DIVIDE(1),
    .CLKOUT5_DUTY_CYCLE(0.5),
    .CLKOUT5_PHASE(0),
    .CLKOUT6_DIVIDE(1),
    .CLKOUT6_DUTY_CYCLE(0.5),
    .CLKOUT6_PHASE(0),
    .CLKFBOUT_MULT_F(5),
    .CLKFBOUT_PHASE(0),
    .DIVCLK_DIVIDE(1),
    .REF_JITTER1(0.010),
    .CLKIN1_PERIOD(5.0),
    .STARTUP_WAIT("FALSE"),
    .CLKOUT4_CASCADE("FALSE")
)
clk_mmcm_inst (
    .CLKIN1(clk_200mhz_ibufg),
    .CLKFBIN(mmcm_clkfb),
    .RST(mmcm_rst),
    .PWRDWN(1'b0),
    .CLKOUT0(clk_mmcm_out),
    .CLKOUT0B(),
    .CLKOUT1(),
    .CLKOUT1B(),
    .CLKOUT2(clk_200mhz_mmcm_out),
    .CLKOUT2B(),
    .CLKOUT3(clk_50mhz_mmcm_out),
    .CLKOUT3B(),
    .CLKOUT4(),
    .CLKOUT5(),
    .CLKOUT6(),
    .CLKFBOUT(mmcm_clkfb),
    .CLKFBOUTB(),
    .LOCKED(mmcm_locked)
);

BUFG
clk_bufg_inst (
    .I(clk_mmcm_out),
    .O(clk_int)
);

// BUFG
// clk_25mhz_bufg_inst (
//     .I(clk_25mhz_mmcm_out),
//     .O(clk_25mhz_int)
// );

BUFG
clk_50mhz_bufg_inst (
    .I(clk_50mhz_mmcm_out),
    .O(clk_50mhz_int)
);

BUFG
clk_200mhz_bufg_inst (
    .I(clk_200mhz_mmcm_out),
    .O(clk_200mhz_int)
);

sync_reset #(
    .N(4)
)
sync_reset_inst (
    .clk(clk_int),
    .rst(~mmcm_locked),
    .out(rst_int)
);

// GPIO
wire btnu_int;
wire btnl_int;
wire btnd_int;
wire btnr_int;
wire btnc_int;
wire [3:0] sw_int;

debounce_switch #(
    .WIDTH(9),
    .N(4),
    .RATE(125000)
)
debounce_switch_inst (
    .clk(clk_int),
    .rst(rst_int),
    .in({btnu,
        btnl,
        btnd,
        btnr,
        btnc,
        sw}),
    .out({btnu_int,
        btnl_int,
        btnd_int,
        btnr_int,
        btnc_int,
        sw_int})
);

wire uart_rxd_int;
wire uart_cts_int;

sync_signal #(
    .WIDTH(2),
    .N(2)
)
sync_signal_inst (
    .clk(clk_int),
    .in({uart_rxd, uart_cts}),
    .out({uart_rxd_int, uart_cts_int})
);

// IODELAY elements for RGMII interface to PHY
// wire [3:0] phy_rxd_delay;
// wire       phy_rx_ctl_delay;

// IDELAYCTRL
// idelayctrl_inst (
//     .REFCLK(clk_200mhz_int),
//     .RST(rst_int),
//     .RDY()
// );

// IDELAYE2 #(
//     .IDELAY_TYPE("FIXED")
// )
// phy_rxd_idelay_0 (
//     .IDATAIN(phy_rxd[0]),
//     .DATAOUT(phy_rxd_delay[0]),
//     .DATAIN(1'b0),
//     .C(1'b0),
//     .CE(1'b0),
//     .INC(1'b0),
//     .CINVCTRL(1'b0),
//     .CNTVALUEIN(5'd0),
//     .CNTVALUEOUT(),
//     .LD(1'b0),
//     .LDPIPEEN(1'b0),
//     .REGRST(1'b0)
// );

// IDELAYE2 #(
//     .IDELAY_TYPE("FIXED")
// )
// phy_rxd_idelay_1 (
//     .IDATAIN(phy_rxd[1]),
//     .DATAOUT(phy_rxd_delay[1]),
//     .DATAIN(1'b0),
//     .C(1'b0),
//     .CE(1'b0),
//     .INC(1'b0),
//     .CINVCTRL(1'b0),
//     .CNTVALUEIN(5'd0),
//     .CNTVALUEOUT(),
//     .LD(1'b0),
//     .LDPIPEEN(1'b0),
//     .REGRST(1'b0)
// );

// IDELAYE2 #(
//     .IDELAY_TYPE("FIXED")
// )
// phy_rxd_idelay_2 (
//     .IDATAIN(phy_rxd[2]),
//     .DATAOUT(phy_rxd_delay[2]),
//     .DATAIN(1'b0),
//     .C(1'b0),
//     .CE(1'b0),
//     .INC(1'b0),
//     .CINVCTRL(1'b0),
//     .CNTVALUEIN(5'd0),
//     .CNTVALUEOUT(),
//     .LD(1'b0),
//     .LDPIPEEN(1'b0),
//     .REGRST(1'b0)
// );

// IDELAYE2 #(
//     .IDELAY_TYPE("FIXED")
// )
// phy_rxd_idelay_3 (
//     .IDATAIN(phy_rxd[3]),
//     .DATAOUT(phy_rxd_delay[3]),
//     .DATAIN(1'b0),
//     .C(1'b0),
//     .CE(1'b0),
//     .INC(1'b0),
//     .CINVCTRL(1'b0),
//     .CNTVALUEIN(5'd0),
//     .CNTVALUEOUT(),
//     .LD(1'b0),
//     .LDPIPEEN(1'b0),
//     .REGRST(1'b0)
// );

// IDELAYE2 #(
//     .IDELAY_TYPE("FIXED")
// )
// phy_rx_ctl_idelay (
//     .IDATAIN(phy_rx_ctl),
//     .DATAOUT(phy_rx_ctl_delay),
//     .DATAIN(1'b0),
//     .C(1'b0),
//     .CE(1'b0),
//     .INC(1'b0),
//     .CINVCTRL(1'b0),
//     .CNTVALUEIN(5'd0),
//     .CNTVALUEOUT(),
//     .LD(1'b0),
//     .LDPIPEEN(1'b0),
//     .REGRST(1'b0)
// );

fpga_core #(
    .TARGET("XILINX")
    //.TARGET("GENERIC")
)
core_inst (
    /*
     * Clock: 125MHz
     * Synchronous reset
     */
    .clk(clk_int),
    .rst(rst_int),
    /*
     * GPIO
     */
    .btnu(btnu_int),
    .btnl(btnl_int),
    .btnd(btnd_int),
    .btnr(btnr_int),
    .btnc(btnc_int),
    .sw(sw_int),
    .led(led_out),
    /*
     * Ethernet: 100BASE-T RMII
     */
    .phy_rxd(phy_rxd),
    .phy_rx_er(phy_rx_er),
    .phy_crs_dv(phy_crs_dv),
    .phy_txd(phy_txd),
    .phy_tx_en(phy_tx_en),
    .phy_ref_clk(clk_50mhz_int),
    .phy_reset_n(phy_reset),
    .phy_int_n(phy_int_n),

    .phy_mii_tx_clk(phy_mii_tx_clk),

    /*
     * UART: 115200 bps, 8N1
     */
    .uart_rxd(uart_rxd_int),
    .uart_txd(uart_txd),
    .uart_rts(uart_rts),
    .uart_cts(uart_cts_int)
);

endmodule

`resetall
